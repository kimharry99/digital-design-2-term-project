module main()
endmodule